
`timescale 1 ps / 1 ps

module system_top(
    DDR_addr,
    DDR_ba,
    DDR_cas_n,
    DDR_ck_n,
    DDR_ck_p,
    DDR_cke,
    DDR_cs_n,
    DDR_dm,
    DDR_dq,
    DDR_dqs_n,
    DDR_dqs_p,
    DDR_odt,
    DDR_ras_n,
    DDR_reset_n,
    DDR_we_n,
    FIXED_IO_ddr_vrn,
    FIXED_IO_ddr_vrp,
    FIXED_IO_mio,
    FIXED_IO_ps_clk,
    FIXED_IO_ps_porb,
    FIXED_IO_ps_srstb,

    GPIO2_0_tri_io,
    GPIO_0_tri_io,
    HDMI_clk_n,
    HDMI_clk_p,
    HDMI_data_n,
    HDMI_data_p,

    led4_b,
    led4_g,
    led4_r,
    led5_b,
    led5_g,
    led5_r
);
    inout [14:0]DDR_addr;
    inout [2:0]DDR_ba;
    inout DDR_cas_n;
    inout DDR_ck_n;
    inout DDR_ck_p;
    inout DDR_cke;
    inout DDR_cs_n;
    inout [3:0]DDR_dm;
    inout [31:0]DDR_dq;
    inout [3:0]DDR_dqs_n;
    inout [3:0]DDR_dqs_p;
    inout DDR_odt;
    inout DDR_ras_n;
    inout DDR_reset_n;
    inout DDR_we_n;
    inout FIXED_IO_ddr_vrn;
    inout FIXED_IO_ddr_vrp;
    inout [53:0]FIXED_IO_mio;
    inout FIXED_IO_ps_clk;
    inout FIXED_IO_ps_porb;
    inout FIXED_IO_ps_srstb;

    inout GPIO2_0_tri_io;
    inout GPIO_0_tri_io;
    output HDMI_clk_n;
    output HDMI_clk_p;
    output [2:0]HDMI_data_n;
    output [2:0]HDMI_data_p;
    output led4_b;
    output led4_g;
    output led4_r;
    output led5_b;
    output led5_g;
    output led5_r;

    wire [14:0]DDR_addr;
    wire [2:0]DDR_ba;
    wire DDR_cas_n;
    wire DDR_ck_n;
    wire DDR_ck_p;
    wire DDR_cke;
    wire DDR_cs_n;
    wire [3:0]DDR_dm;
    wire [31:0]DDR_dq;
    wire [3:0]DDR_dqs_n;
    wire [3:0]DDR_dqs_p;
    wire DDR_odt;
    wire DDR_ras_n;
    wire DDR_reset_n;
    wire DDR_we_n;
    wire FIXED_IO_ddr_vrn;
    wire FIXED_IO_ddr_vrp;
    wire [53:0]FIXED_IO_mio;
    wire FIXED_IO_ps_clk;
    wire FIXED_IO_ps_porb;
    wire FIXED_IO_ps_srstb;

    wire GPIO2_0_tri_io;
    wire GPIO_0_tri_io;
    wire HDMI_clk_n;
    wire HDMI_clk_p;
    wire [2:0]HDMI_data_n;
    wire [2:0]HDMI_data_p;
    wire [5:0]rgb;

    assign 
        led4_b = rgb[5],
        led4_g = rgb[4],
        led4_r = rgb[3],
        led5_b = rgb[2],
        led5_g = rgb[1],
        led5_r = rgb[0];
    
    system_wrapper i_system_wrapper (
        .DDR_addr(DDR_addr),
        .DDR_ba(DDR_ba),
        .DDR_cas_n(DDR_cas_n),
        .DDR_ck_n(DDR_ck_n),
        .DDR_ck_p(DDR_ck_p),
        .DDR_cke(DDR_cke),
        .DDR_cs_n(DDR_cs_n),
        .DDR_dm(DDR_dm),
        .DDR_dq(DDR_dq),
        .DDR_dqs_n(DDR_dqs_n),
        .DDR_dqs_p(DDR_dqs_p),
        .DDR_odt(DDR_odt),
        .DDR_ras_n(DDR_ras_n),
        .DDR_reset_n(DDR_reset_n),
        .DDR_we_n(DDR_we_n),
        .FIXED_IO_ddr_vrn(FIXED_IO_ddr_vrn),
        .FIXED_IO_ddr_vrp(FIXED_IO_ddr_vrp),
        .FIXED_IO_mio(FIXED_IO_mio),
        .FIXED_IO_ps_clk(FIXED_IO_ps_clk),
        .FIXED_IO_ps_porb(FIXED_IO_ps_porb),
        .FIXED_IO_ps_srstb(FIXED_IO_ps_srstb),
        .GPIO2_0_tri_io(GPIO2_0_tri_io),
        .GPIO_0_tri_io(GPIO_0_tri_io),
        .HDMI_clk_n(HDMI_clk_n),
        .HDMI_clk_p(HDMI_clk_p),
        .HDMI_data_n(HDMI_data_n),
        .HDMI_data_p(HDMI_data_p),
        .rgb(rgb)
    );

endmodule
