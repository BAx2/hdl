`ifndef CORDIC_SVH
`define CORDIC_SVH

parameter CORDIC_SCALE_K = 1.64676026;

`endif